module stripe(
	      
	      );
endmodule // stripe
