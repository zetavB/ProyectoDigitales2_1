module serial_parallel(

);

endmodule