module conv8_32(
		
		);
endmodule // conv8_32
