module unstripe(
		
		);
endmodule // unstripe
