module genClock(
		
		);
endmodule // genClock
