module conv32_8(
		
		);
endmodule // conv32_8
